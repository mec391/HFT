module hft(

input clk,
input rx,
output tx

	);

reset_n = 1'b1;


//instantiate the UART modules
uart uu0(


	);

//instantiate the addr mux

//instantiate the system addr 0
		//FOR ADDR 0:
		//instantiate DP-BRAM (Book Handler)
		//instantiate MA algo
		//instantiate NN1 algo
		//instantiate NN2 algo
		//instantiate decision-making module
		//instantiate timestamp

endmodule

