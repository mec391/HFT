module tx_mux(


);


endmodule