module timestamp(


);


endmodule