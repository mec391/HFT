module ema(



);





endmodule


module four_sec_timer(
input clk,
input reset_n,
output reg sec_dv
	);




endmodule

module bid_ask_averager(



	);


endmodule